��m o d u l e   b r a u n _ m u l t i p l i e r _ t b _ t o p ;  
         l o g i c   [ 1 : 0 ]   a ,   b ;  
         o u t p u t   [ 2 : 0 ]   p ;  
          
         b r a u n _ m u l t i p l i e r   d u t   ( a ,   b ,   p ) ;  
  
         i n i t i a l   b e g i n  
                 / /   T e s t   c a s e   1 :   0   *   0   =   0  
                 a   =   2 ' b 0 0 ;   b   =   2 ' b 0 0 ;  
                 # 1 0 ;  
                 a s s e r t   ( p   = =   3 ' b 0 0 0 )   e l s e   $ f a t a l ( " T e s t   c a s e   1   f a i l e d :   % b   *   % b   =   % b " ,   a ,   b ,   p ) ;  
  
                 / /   T e s t   c a s e   2 :   0   *   1   =   0  
                 a   =   2 ' b 0 0 ;   b   =   2 ' b 0 1 ;  
                 # 1 0 ;  
                 a s s e r t   ( p   = =   3 ' b 0 0 0 )   e l s e   $ f a t a l ( " T e s t   c a s e   2   f a i l e d :   % b   *   % b   =   % b " ,   a ,   b ,   p ) ;  
  
                 / /   T e s t   c a s e   3 :   1   *   0   =   0  
                 a   =   2 ' b 0 1 ;   b   =   2 ' b 0 0 ;  
                 # 1 0 ;  
                 a s s e r t   ( p   = =   3 ' b 0 0 0 )   e l s e   $ f a t a l ( " T e s t   c a s e   3   f a i l e d :   % b   *   % b   =   % b " ,   a ,   b ,   p ) ;  
  
                 / /   T e s t   c a s e   4 :   1   *   1   =   1  
                 a   =   2 ' b 0 1 ;   b   =   2 ' b 0 1 ;  
                 # 1 0 ;  
                 a s s e r t   ( p   = =   3 ' b 0 0 1 )   e l s e   $ f a t a l ( " T e s t   c a s e   4   f a i l e d :   % b   *   % b   =   % b " ,   a ,   b ,   p ) ;  
  
                 / /   T e s t   c a s e   5 :   1   *   2   =   2  
                 a   =   2 ' b 0 1 ;   b   =   2 ' b 1 0 ;  
                 # 1 0 ;  
                 a s s e r t   ( p   = =   3 ' b 0 1 0 )   e l s e   $ f a t a l ( " T e s t   c a s e   5   f a i l e d :   % b   *   % b   =   % b " ,   a ,   b ,   p ) ;  
  
                 / /   T e s t   c a s e   6 :   2   *   1   =   2  
                 a   =   2 ' b 1 0 ;   b   =   2 ' b 0 1 ;  
                 # 1 0 ;  
                 a s s e r t   ( p   = =   3 ' b 0 1 0 )   e l s e   $ f a t a l ( " T e s t   c a s e   6   f a i l e d :   % b   *   % b   =   % b " ,   a ,   b ,   p ) ;  
  
                 / /   T e s t   c a s e   7 :   M a x   v a l u e   t e s t :   ( 3 * 3 = 9 )  
                 a   =   ' h 1 1 ;   b   =   ' h 1 1 ;  
                 # 1 0 ;  
                 a s s e r t   ( p   = =   ' h 1 0 0 1 )   e l s e   $ f a t a l ( " T e s t   c a s e   m a x   v a l u e   f a i l e d :   % h   *   % h   ! =   % h " ,   a ,   b ,   p ) ;  
                  
         e n d  
 e n d m o d u l e 